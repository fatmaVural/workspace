//Design and simulate  a decoder for  7 segment display.

module display7seg_main(A,Y);

input [3:0] A;
output [6:0] Y;

wire [3:0] A;
wire [6:0] Y;

assign Y[6] = (~A[3] & ~A[2] & ~A[1] & ~A[0]) | (~A[3] & ~A[2] & ~A[1] & A[0])| 
            (~A[3] & A[2] & A[1] & A[0])|(A[3] & A[2] & ~A[1] & ~A[0]);
				
assign Y[5]=(~A[3] & ~A[2] & ~A[1] & A[0]) | (~A[3] & ~A[2] & A[1] & ~A[0])| 
            (~A[3] & ~A[2] & A[1] & A[0])|(~A[3] & A[2] & A[1] & A[0])|(A[3] & A[2] & ~A[1] & A[0]);
	
assign Y[4]=(~A[3] & ~A[2] & ~A[1] & A[0]) | (~A[3] & ~A[2] & A[1] & A[0]) | 
            (~A[3] & A[2] & ~A[1] & ~A[0]) | (~A[3] & A[2] & ~A[1] & A[0]) | 
				(~A[3] & A[2] & A[1] & A[0]) | (A[3] & ~A[2] & ~A[1] & A[0]);
				
assign Y[3]=(~A[3] & ~A[2] & ~A[1] & A[0]) | (~A[3] & A[2] & ~A[1] & ~A[0])| 
            (~A[3] & A[2] & A[1] & A[0])|(A[3] & ~A[2] & ~A[1] & A[0]) |(A[3] & ~A[2] & A[1] & ~A[0])|
				(A[3] & A[2] & A[1] & A[0]);
			

assign Y[2]=(~A[3] & ~A[2] & A[1] & ~A[0]) | (A[3] & A[2] & ~A[1] & ~A[0])| 
            (A[3] & A[2] & A[1] & ~A[0]) | (A[3] & A[2] & A[1] & A[0]);
				
//assign Y[1]=(~A[3] & A[2] & ~A[1] & A[0]) | (A[3] & A[2] & ~A[1] & ~A[0])| (A[3] &  A[1] & A[0])|(A[2] & A[1] & ~A[0]);
assign Y[1]= (~A[3] & A[2] & ~A[1] & A[0]) | (~A[3] & A[2] & A[1] & ~A[0])| 
            (A[3] & ~A[2] & A[1] & A[0])|(A[3] & A[2] & ~A[1] & ~A[0]) | (A[3] & A[2] & A[1] & ~A[0]) |
				(A[3] & A[2] & A[1] & A[0]);

				
assign Y[0]=(~A[3] & ~A[2] & ~A[1] & A[0]) | (~A[3] & A[2] & ~A[1] & ~A[0])| 
            (A[3] & ~A[2] & A[1] & A[0]) | (A[3] & A[2] & ~A[1] & A[0]);
				
endmodule
