library verilog;
use verilog.vl_types.all;
entity johnson_8bit_tb is
    generic(
        period          : integer := 20
    );
end johnson_8bit_tb;
