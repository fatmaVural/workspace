library verilog;
use verilog.vl_types.all;
entity lpm_shiftreg0_tb is
    generic(
        period          : integer := 20
    );
end lpm_shiftreg0_tb;
