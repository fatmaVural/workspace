//testbench
`timescale 1ns/1ps
module comperator_testbench();

reg [7:0]A;
reg [7:0]B;
wire C,D;

comperator_main UUt(.A(A),.B(B),.C(C),.D(D));

initial
begin
A <= 8'b00000001; 
B <= 8'b00000000; #10;
A <= 8'b00000010; #10;
B <= 8'b00000010; #10;
A <= 8'b00000110; #10;
B <= 8'b00000010; #10;
A <= 8'b00000101; #10;
B <= 8'b00000010; #10;
A <= 8'b10101010; #10;
B <= 8'b11111101; #10;
A <= 8'b11111101; #10;
B <= 8'b10000010; #10;
A <= 8'b11000000; #10;
B <= 8'b00001110; #10;
A <= 8'b11000000; #10;
B <= 8'b11111111; #10;
A <= 8'b11111110; #10;
B <= 8'b11111111; #10;
end
endmodule 
